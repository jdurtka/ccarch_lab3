library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


--LUT concept derived from http://stackoverflow.com/questions/21976749/design-of-a-vhdl-lut-module

--Implements an 8 bit x 32 bit LUT (truncates input and output fractions accordingly)

--Values generated using the Matlab script LUT_gen.m

entity LUT is
    port (
			clk : in std_logic;
			x_beta : in std_logic_vector(27 downto 0);
			x_beta_lut_out : out std_logic_vector(27 downto 0)
    );

	constant W : integer := 28;
	constant F : integer := 14;

end entity;

architecture LUT_arch of LUT is
	signal x_beta_part : std_logic_vector(13 downto 6);
	signal x_beta_lut : std_logic_vector(31 downto 0);
begin

		x_beta_part <= x_beta(13 downto 6);
		x_beta_lut_out <= x_beta_lut(31 downto 4);

    process (clk) is
    begin
			if (rising_edge(clk)) then
        case (x_beta_part) is      
			--when "0000" => xyz <= "000" ;
			-- 1.000000 => 1.000000
			when "00000000" => x_beta_lut <= "00000000000001000000000000000000" ;
			-- 1.003906 => 0.994167
			when "00000001" => x_beta_lut <= "00000000000000111111101000000111" ;
			-- 1.007813 => 0.988396
			when "00000010" => x_beta_lut <= "00000000000000111111010000011110" ;
			-- 1.011719 => 0.982677
			when "00000011" => x_beta_lut <= "00000000000000111110111001000011" ;
			-- 1.015625 => 0.977013
			when "00000100" => x_beta_lut <= "00000000000000111110100001110110" ;
			-- 1.019531 => 0.971401
			when "00000101" => x_beta_lut <= "00000000000000111110001010110111" ;
			-- 1.023438 => 0.965847
			when "00000110" => x_beta_lut <= "00000000000000111101110100000111" ;
			-- 1.027344 => 0.960342
			when "00000111" => x_beta_lut <= "00000000000000111101011101100100" ;
			-- 1.031250 => 0.954891
			when "00001000" => x_beta_lut <= "00000000000000111101000111001111" ;
			-- 1.035156 => 0.949493
			when "00001001" => x_beta_lut <= "00000000000000111100110001001000" ;
			-- 1.039063 => 0.944141
			when "00001010" => x_beta_lut <= "00000000000000111100011011001101" ;
			-- 1.042969 => 0.938843
			when "00001011" => x_beta_lut <= "00000000000000111100000101100000" ;
			-- 1.046875 => 0.933594
			when "00001100" => x_beta_lut <= "00000000000000111011110000000000" ;
			-- 1.050781 => 0.928391
			when "00001101" => x_beta_lut <= "00000000000000111011011010101100" ;
			-- 1.054688 => 0.923241
			when "00001110" => x_beta_lut <= "00000000000000111011000101100110" ;
			-- 1.058594 => 0.918133
			when "00001111" => x_beta_lut <= "00000000000000111010110000101011" ;
			-- 1.062500 => 0.913074
			when "00010000" => x_beta_lut <= "00000000000000111010011011111101" ;
			-- 1.066406 => 0.908062
			when "00010001" => x_beta_lut <= "00000000000000111010000111011011" ;
			-- 1.070313 => 0.903095
			when "00010010" => x_beta_lut <= "00000000000000111001110011000101" ;
			-- 1.074219 => 0.898174
			when "00010011" => x_beta_lut <= "00000000000000111001011110111011" ;
			-- 1.078125 => 0.893299
			when "00010100" => x_beta_lut <= "00000000000000111001001010111101" ;
			-- 1.082031 => 0.888466
			when "00010101" => x_beta_lut <= "00000000000000111000110111001010" ;
			-- 1.085938 => 0.883675
			when "00010110" => x_beta_lut <= "00000000000000111000100011100010" ;
			-- 1.089844 => 0.878929
			when "00010111" => x_beta_lut <= "00000000000000111000010000000110" ;
			-- 1.093750 => 0.874226
			when "00011000" => x_beta_lut <= "00000000000000110111111100110101" ;
			-- 1.097656 => 0.869560
			when "00011001" => x_beta_lut <= "00000000000000110111101001101110" ;
			-- 1.101563 => 0.864941
			when "00011010" => x_beta_lut <= "00000000000000110111010110110011" ;
			-- 1.105469 => 0.860359
			when "00011011" => x_beta_lut <= "00000000000000110111000100000010" ;
			-- 1.109375 => 0.855820
			when "00011100" => x_beta_lut <= "00000000000000110110110001011100" ;
			-- 1.113281 => 0.851318
			when "00011101" => x_beta_lut <= "00000000000000110110011111000000" ;
			-- 1.117188 => 0.846859
			when "00011110" => x_beta_lut <= "00000000000000110110001100101111" ;
			-- 1.121094 => 0.842438
			when "00011111" => x_beta_lut <= "00000000000000110101111010101000" ;
			-- 1.125000 => 0.838051
			when "00100000" => x_beta_lut <= "00000000000000110101101000101010" ;
			-- 1.128906 => 0.833706
			when "00100001" => x_beta_lut <= "00000000000000110101010110110111" ;
			-- 1.132813 => 0.829399
			when "00100010" => x_beta_lut <= "00000000000000110101000101001110" ;
			-- 1.136719 => 0.825127
			when "00100011" => x_beta_lut <= "00000000000000110100110011101110" ;
			-- 1.140625 => 0.820892
			when "00100100" => x_beta_lut <= "00000000000000110100100010011000" ;
			-- 1.144531 => 0.816692
			when "00100101" => x_beta_lut <= "00000000000000110100010001001011" ;
			-- 1.148438 => 0.812531
			when "00100110" => x_beta_lut <= "00000000000000110100000000001000" ;
			-- 1.152344 => 0.808403
			when "00100111" => x_beta_lut <= "00000000000000110011101111001110" ;
			-- 1.156250 => 0.804310
			when "00101000" => x_beta_lut <= "00000000000000110011011110011101" ;
			-- 1.160156 => 0.800251
			when "00101001" => x_beta_lut <= "00000000000000110011001101110101" ;
			-- 1.164063 => 0.796223
			when "00101010" => x_beta_lut <= "00000000000000110010111101010101" ;
			-- 1.167969 => 0.792233
			when "00101011" => x_beta_lut <= "00000000000000110010101100111111" ;
			-- 1.171875 => 0.788277
			when "00101100" => x_beta_lut <= "00000000000000110010011100110010" ;
			-- 1.175781 => 0.784351
			when "00101101" => x_beta_lut <= "00000000000000110010001100101101" ;
			-- 1.179688 => 0.780457
			when "00101110" => x_beta_lut <= "00000000000000110001111100110000" ;
			-- 1.183594 => 0.776596
			when "00101111" => x_beta_lut <= "00000000000000110001101100111100" ;
			-- 1.187500 => 0.772770
			when "00110000" => x_beta_lut <= "00000000000000110001011101010001" ;
			-- 1.191406 => 0.768970
			when "00110001" => x_beta_lut <= "00000000000000110001001101101101" ;
			-- 1.195313 => 0.765205
			when "00110010" => x_beta_lut <= "00000000000000110000111110010010" ;
			-- 1.199219 => 0.761471
			when "00110011" => x_beta_lut <= "00000000000000110000101110111111" ;
			-- 1.203125 => 0.757763
			when "00110100" => x_beta_lut <= "00000000000000110000011111110011" ;
			-- 1.207031 => 0.754089
			when "00110101" => x_beta_lut <= "00000000000000110000010000110000" ;
			-- 1.210938 => 0.750443
			when "00110110" => x_beta_lut <= "00000000000000110000000001110100" ;
			-- 1.214844 => 0.746826
			when "00110111" => x_beta_lut <= "00000000000000101111110011000000" ;
			-- 1.218750 => 0.743237
			when "00111000" => x_beta_lut <= "00000000000000101111100100010011" ;
			-- 1.222656 => 0.739677
			when "00111001" => x_beta_lut <= "00000000000000101111010101101110" ;
			-- 1.226563 => 0.736149
			when "00111010" => x_beta_lut <= "00000000000000101111000111010001" ;
			-- 1.230469 => 0.732647
			when "00111011" => x_beta_lut <= "00000000000000101110111000111011" ;
			-- 1.234375 => 0.729172
			when "00111100" => x_beta_lut <= "00000000000000101110101010101100" ;
			-- 1.238281 => 0.725723
			when "00111101" => x_beta_lut <= "00000000000000101110011100100100" ;
			-- 1.242188 => 0.722301
			when "00111110" => x_beta_lut <= "00000000000000101110001110100011" ;
			-- 1.246094 => 0.718910
			when "00111111" => x_beta_lut <= "00000000000000101110000000101010" ;
			-- 1.250000 => 0.715542
			when "01000000" => x_beta_lut <= "00000000000000101101110010110111" ;
			-- 1.253906 => 0.712200
			when "01000001" => x_beta_lut <= "00000000000000101101100101001011" ;
			-- 1.257813 => 0.708885
			when "01000010" => x_beta_lut <= "00000000000000101101010111100110" ;
			-- 1.261719 => 0.705597
			when "01000011" => x_beta_lut <= "00000000000000101101001010001000" ;
			-- 1.265625 => 0.702332
			when "01000100" => x_beta_lut <= "00000000000000101100111100110000" ;
			-- 1.269531 => 0.699093
			when "01000101" => x_beta_lut <= "00000000000000101100101111011111" ;
			-- 1.273438 => 0.695877
			when "01000110" => x_beta_lut <= "00000000000000101100100010010100" ;
			-- 1.277344 => 0.692688
			when "01000111" => x_beta_lut <= "00000000000000101100010101010000" ;
			-- 1.281250 => 0.689522
			when "01001000" => x_beta_lut <= "00000000000000101100001000010010" ;
			-- 1.285156 => 0.686382
			when "01001001" => x_beta_lut <= "00000000000000101011111011011011" ;
			-- 1.289063 => 0.683266
			when "01001010" => x_beta_lut <= "00000000000000101011101110101010" ;
			-- 1.292969 => 0.680172
			when "01001011" => x_beta_lut <= "00000000000000101011100001111111" ;
			-- 1.296875 => 0.677101
			when "01001100" => x_beta_lut <= "00000000000000101011010101011010" ;
			-- 1.300781 => 0.674053
			when "01001101" => x_beta_lut <= "00000000000000101011001000111011" ;
			-- 1.304688 => 0.671028
			when "01001110" => x_beta_lut <= "00000000000000101010111100100010" ;
			-- 1.308594 => 0.668026
			when "01001111" => x_beta_lut <= "00000000000000101010110000001111" ;
			-- 1.312500 => 0.665047
			when "01010000" => x_beta_lut <= "00000000000000101010100100000010" ;
			-- 1.316406 => 0.662086
			when "01010001" => x_beta_lut <= "00000000000000101010010111111010" ;
			-- 1.320313 => 0.659149
			when "01010010" => x_beta_lut <= "00000000000000101010001011111000" ;
			-- 1.324219 => 0.656235
			when "01010011" => x_beta_lut <= "00000000000000101001111111111100" ;
			-- 1.328125 => 0.653343
			when "01010100" => x_beta_lut <= "00000000000000101001110100000110" ;
			-- 1.332031 => 0.650471
			when "01010101" => x_beta_lut <= "00000000000000101001101000010101" ;
			-- 1.335938 => 0.647621
			when "01010110" => x_beta_lut <= "00000000000000101001011100101010" ;
			-- 1.339844 => 0.644791
			when "01010111" => x_beta_lut <= "00000000000000101001010001000100" ;
			-- 1.343750 => 0.641983
			when "01011000" => x_beta_lut <= "00000000000000101001000101100100" ;
			-- 1.347656 => 0.639191
			when "01011001" => x_beta_lut <= "00000000000000101000111010001000" ;
			-- 1.351563 => 0.636421
			when "01011010" => x_beta_lut <= "00000000000000101000101110110010" ;
			-- 1.355469 => 0.633675
			when "01011011" => x_beta_lut <= "00000000000000101000100011100010" ;
			-- 1.359375 => 0.630943
			when "01011100" => x_beta_lut <= "00000000000000101000011000010110" ;
			-- 1.363281 => 0.628235
			when "01011101" => x_beta_lut <= "00000000000000101000001101010000" ;
			-- 1.367188 => 0.625546
			when "01011110" => x_beta_lut <= "00000000000000101000000010001111" ;
			-- 1.371094 => 0.622871
			when "01011111" => x_beta_lut <= "00000000000000100111110111010010" ;
			-- 1.375000 => 0.620220
			when "01100000" => x_beta_lut <= "00000000000000100111101100011011" ;
			-- 1.378906 => 0.617588
			when "01100001" => x_beta_lut <= "00000000000000100111100001101001" ;
			-- 1.382813 => 0.614971
			when "01100010" => x_beta_lut <= "00000000000000100111010110111011" ;
			-- 1.386719 => 0.612373
			when "01100011" => x_beta_lut <= "00000000000000100111001100010010" ;
			-- 1.390625 => 0.609798
			when "01100100" => x_beta_lut <= "00000000000000100111000001101111" ;
			-- 1.394531 => 0.607235
			when "01100101" => x_beta_lut <= "00000000000000100110110111001111" ;
			-- 1.398438 => 0.604694
			when "01100110" => x_beta_lut <= "00000000000000100110101100110101" ;
			-- 1.402344 => 0.602169
			when "01100111" => x_beta_lut <= "00000000000000100110100010011111" ;
			-- 1.406250 => 0.599663
			when "01101000" => x_beta_lut <= "00000000000000100110011000001110" ;
			-- 1.410156 => 0.597172
			when "01101001" => x_beta_lut <= "00000000000000100110001110000001" ;
			-- 1.414063 => 0.594700
			when "01101010" => x_beta_lut <= "00000000000000100110000011111001" ;
			-- 1.417969 => 0.592243
			when "01101011" => x_beta_lut <= "00000000000000100101111001110101" ;
			-- 1.421875 => 0.589806
			when "01101100" => x_beta_lut <= "00000000000000100101101111110110" ;
			-- 1.425781 => 0.587383
			when "01101101" => x_beta_lut <= "00000000000000100101100101111011" ;
			-- 1.429688 => 0.584976
			when "01101110" => x_beta_lut <= "00000000000000100101011100000100" ;
			-- 1.433594 => 0.582588
			when "01101111" => x_beta_lut <= "00000000000000100101010010010010" ;
			-- 1.437500 => 0.580215
			when "01110000" => x_beta_lut <= "00000000000000100101001000100100" ;
			-- 1.441406 => 0.577858
			when "01110001" => x_beta_lut <= "00000000000000100100111110111010" ;
			-- 1.445313 => 0.575516
			when "01110010" => x_beta_lut <= "00000000000000100100110101010100" ;
			-- 1.449219 => 0.573189
			when "01110011" => x_beta_lut <= "00000000000000100100101011110010" ;
			-- 1.453125 => 0.570881
			when "01110100" => x_beta_lut <= "00000000000000100100100010010101" ;
			-- 1.457031 => 0.568588
			when "01110101" => x_beta_lut <= "00000000000000100100011000111100" ;
			-- 1.460938 => 0.566307
			when "01110110" => x_beta_lut <= "00000000000000100100001111100110" ;
			-- 1.464844 => 0.564045
			when "01110111" => x_beta_lut <= "00000000000000100100000110010101" ;
			-- 1.468750 => 0.561794
			when "01111000" => x_beta_lut <= "00000000000000100011111101000111" ;
			-- 1.472656 => 0.559563
			when "01111001" => x_beta_lut <= "00000000000000100011110011111110" ;
			-- 1.476563 => 0.557343
			when "01111010" => x_beta_lut <= "00000000000000100011101010111000" ;
			-- 1.480469 => 0.555138
			when "01111011" => x_beta_lut <= "00000000000000100011100001110110" ;
			-- 1.484375 => 0.552948
			when "01111100" => x_beta_lut <= "00000000000000100011011000111000" ;
			-- 1.488281 => 0.550774
			when "01111101" => x_beta_lut <= "00000000000000100011001111111110" ;
			-- 1.492188 => 0.548611
			when "01111110" => x_beta_lut <= "00000000000000100011000111000111" ;
			-- 1.496094 => 0.546463
			when "01111111" => x_beta_lut <= "00000000000000100010111110010100" ;
			-- 1.500000 => 0.544331
			when "10000000" => x_beta_lut <= "00000000000000100010110101100101" ;
			-- 1.503906 => 0.542213
			when "10000001" => x_beta_lut <= "00000000000000100010101100111010" ;
			-- 1.507813 => 0.540108
			when "10000010" => x_beta_lut <= "00000000000000100010100100010010" ;
			-- 1.511719 => 0.538013
			when "10000011" => x_beta_lut <= "00000000000000100010011011101101" ;
			-- 1.515625 => 0.535934
			when "10000100" => x_beta_lut <= "00000000000000100010010011001100" ;
			-- 1.519531 => 0.533871
			when "10000101" => x_beta_lut <= "00000000000000100010001010101111" ;
			-- 1.523438 => 0.531818
			when "10000110" => x_beta_lut <= "00000000000000100010000010010101" ;
			-- 1.527344 => 0.529778
			when "10000111" => x_beta_lut <= "00000000000000100001111001111110" ;
			-- 1.531250 => 0.527752
			when "10001000" => x_beta_lut <= "00000000000000100001110001101011" ;
			-- 1.535156 => 0.525742
			when "10001001" => x_beta_lut <= "00000000000000100001101001011100" ;
			-- 1.539063 => 0.523739
			when "10001010" => x_beta_lut <= "00000000000000100001100001001111" ;
			-- 1.542969 => 0.521751
			when "10001011" => x_beta_lut <= "00000000000000100001011001000110" ;
			-- 1.546875 => 0.519775
			when "10001100" => x_beta_lut <= "00000000000000100001010001000000" ;
			-- 1.550781 => 0.517815
			when "10001101" => x_beta_lut <= "00000000000000100001001000111110" ;
			-- 1.554688 => 0.515865
			when "10001110" => x_beta_lut <= "00000000000000100001000000111111" ;
			-- 1.558594 => 0.513927
			when "10001111" => x_beta_lut <= "00000000000000100000111001000011" ;
			-- 1.562500 => 0.512001
			when "10010000" => x_beta_lut <= "00000000000000100000110001001010" ;
			-- 1.566406 => 0.510086
			when "10010001" => x_beta_lut <= "00000000000000100000101001010100" ;
			-- 1.570313 => 0.508183
			when "10010010" => x_beta_lut <= "00000000000000100000100001100001" ;
			-- 1.574219 => 0.506294
			when "10010011" => x_beta_lut <= "00000000000000100000011001110010" ;
			-- 1.578125 => 0.504414
			when "10010100" => x_beta_lut <= "00000000000000100000010010000101" ;
			-- 1.582031 => 0.502548
			when "10010101" => x_beta_lut <= "00000000000000100000001010011100" ;
			-- 1.585938 => 0.500690
			when "10010110" => x_beta_lut <= "00000000000000100000000010110101" ;
			-- 1.589844 => 0.498848
			when "10010111" => x_beta_lut <= "00000000000000011111111011010010" ;
			-- 1.593750 => 0.497017
			when "10011000" => x_beta_lut <= "00000000000000011111110011110010" ;
			-- 1.597656 => 0.495193
			when "10011001" => x_beta_lut <= "00000000000000011111101100010100" ;
			-- 1.601563 => 0.493382
			when "10011010" => x_beta_lut <= "00000000000000011111100100111001" ;
			-- 1.605469 => 0.491585
			when "10011011" => x_beta_lut <= "00000000000000011111011101100010" ;
			-- 1.609375 => 0.489796
			when "10011100" => x_beta_lut <= "00000000000000011111010110001101" ;
			-- 1.613281 => 0.488018
			when "10011101" => x_beta_lut <= "00000000000000011111001110111011" ;
			-- 1.617188 => 0.486248
			when "10011110" => x_beta_lut <= "00000000000000011111000111101011" ;
			-- 1.621094 => 0.484493
			when "10011111" => x_beta_lut <= "00000000000000011111000000011111" ;
			-- 1.625000 => 0.482746
			when "10100000" => x_beta_lut <= "00000000000000011110111001010101" ;
			-- 1.628906 => 0.481010
			when "10100001" => x_beta_lut <= "00000000000000011110110010001110" ;
			-- 1.632813 => 0.479286
			when "10100010" => x_beta_lut <= "00000000000000011110101011001010" ;
			-- 1.636719 => 0.477573
			when "10100011" => x_beta_lut <= "00000000000000011110100100001001" ;
			-- 1.640625 => 0.475868
			when "10100100" => x_beta_lut <= "00000000000000011110011101001010" ;
			-- 1.644531 => 0.474174
			when "10100101" => x_beta_lut <= "00000000000000011110010110001110" ;
			-- 1.648438 => 0.472488
			when "10100110" => x_beta_lut <= "00000000000000011110001111010100" ;
			-- 1.652344 => 0.470814
			when "10100111" => x_beta_lut <= "00000000000000011110001000011101" ;
			-- 1.656250 => 0.469151
			when "10101000" => x_beta_lut <= "00000000000000011110000001101001" ;
			-- 1.660156 => 0.467495
			when "10101001" => x_beta_lut <= "00000000000000011101111010110111" ;
			-- 1.664063 => 0.465851
			when "10101010" => x_beta_lut <= "00000000000000011101110100001000" ;
			-- 1.667969 => 0.464214
			when "10101011" => x_beta_lut <= "00000000000000011101101101011011" ;
			-- 1.671875 => 0.462589
			when "10101100" => x_beta_lut <= "00000000000000011101100110110001" ;
			-- 1.675781 => 0.460972
			when "10101101" => x_beta_lut <= "00000000000000011101100000001001" ;
			-- 1.679688 => 0.459366
			when "10101110" => x_beta_lut <= "00000000000000011101011001100100" ;
			-- 1.683594 => 0.457767
			when "10101111" => x_beta_lut <= "00000000000000011101010011000001" ;
			-- 1.687500 => 0.456177
			when "10110000" => x_beta_lut <= "00000000000000011101001100100000" ;
			-- 1.691406 => 0.454597
			when "10110001" => x_beta_lut <= "00000000000000011101000110000010" ;
			-- 1.695313 => 0.453030
			when "10110010" => x_beta_lut <= "00000000000000011100111111100111" ;
			-- 1.699219 => 0.451466
			when "10110011" => x_beta_lut <= "00000000000000011100111001001101" ;
			-- 1.703125 => 0.449913
			when "10110100" => x_beta_lut <= "00000000000000011100110010110110" ;
			-- 1.707031 => 0.448372
			when "10110101" => x_beta_lut <= "00000000000000011100101100100010" ;
			-- 1.710938 => 0.446838
			when "10110110" => x_beta_lut <= "00000000000000011100100110010000" ;
			-- 1.714844 => 0.445313
			when "10110111" => x_beta_lut <= "00000000000000011100100000000000" ;
			-- 1.718750 => 0.443794
			when "10111000" => x_beta_lut <= "00000000000000011100011001110010" ;
			-- 1.722656 => 0.442284
			when "10111001" => x_beta_lut <= "00000000000000011100010011100110" ;
			-- 1.726563 => 0.440784
			when "10111010" => x_beta_lut <= "00000000000000011100001101011101" ;
			-- 1.730469 => 0.439293
			when "10111011" => x_beta_lut <= "00000000000000011100000111010110" ;
			-- 1.734375 => 0.437809
			when "10111100" => x_beta_lut <= "00000000000000011100000001010001" ;
			-- 1.738281 => 0.436337
			when "10111101" => x_beta_lut <= "00000000000000011011111011001111" ;
			-- 1.742188 => 0.434868
			when "10111110" => x_beta_lut <= "00000000000000011011110101001110" ;
			-- 1.746094 => 0.433411
			when "10111111" => x_beta_lut <= "00000000000000011011101111010000" ;
			-- 1.750000 => 0.431961
			when "11000000" => x_beta_lut <= "00000000000000011011101001010100" ;
			-- 1.753906 => 0.430515
			when "11000001" => x_beta_lut <= "00000000000000011011100011011001" ;
			-- 1.757813 => 0.429081
			when "11000010" => x_beta_lut <= "00000000000000011011011101100001" ;
			-- 1.761719 => 0.427658
			when "11000011" => x_beta_lut <= "00000000000000011011010111101100" ;
			-- 1.765625 => 0.426239
			when "11000100" => x_beta_lut <= "00000000000000011011010001111000" ;
			-- 1.769531 => 0.424828
			when "11000101" => x_beta_lut <= "00000000000000011011001100000110" ;
			-- 1.773438 => 0.423424
			when "11000110" => x_beta_lut <= "00000000000000011011000110010110" ;
			-- 1.777344 => 0.422031
			when "11000111" => x_beta_lut <= "00000000000000011011000000101001" ;
			-- 1.781250 => 0.420643
			when "11001000" => x_beta_lut <= "00000000000000011010111010111101" ;
			-- 1.785156 => 0.419262
			when "11001001" => x_beta_lut <= "00000000000000011010110101010011" ;
			-- 1.789063 => 0.417889
			when "11001010" => x_beta_lut <= "00000000000000011010101111101011" ;
			-- 1.792969 => 0.416523
			when "11001011" => x_beta_lut <= "00000000000000011010101010000101" ;
			-- 1.796875 => 0.415169
			when "11001100" => x_beta_lut <= "00000000000000011010100100100010" ;
			-- 1.800781 => 0.413818
			when "11001101" => x_beta_lut <= "00000000000000011010011111000000" ;
			-- 1.804688 => 0.412476
			when "11001110" => x_beta_lut <= "00000000000000011010011001100000" ;
			-- 1.808594 => 0.411140
			when "11001111" => x_beta_lut <= "00000000000000011010010100000010" ;
			-- 1.812500 => 0.409809
			when "11010000" => x_beta_lut <= "00000000000000011010001110100101" ;
			-- 1.816406 => 0.408489
			when "11010001" => x_beta_lut <= "00000000000000011010001001001011" ;
			-- 1.820313 => 0.407173
			when "11010010" => x_beta_lut <= "00000000000000011010000011110010" ;
			-- 1.824219 => 0.405869
			when "11010011" => x_beta_lut <= "00000000000000011001111110011100" ;
			-- 1.828125 => 0.404568
			when "11010100" => x_beta_lut <= "00000000000000011001111001000111" ;
			-- 1.832031 => 0.403275
			when "11010101" => x_beta_lut <= "00000000000000011001110011110100" ;
			-- 1.835938 => 0.401989
			when "11010110" => x_beta_lut <= "00000000000000011001101110100011" ;
			-- 1.839844 => 0.400707
			when "11010111" => x_beta_lut <= "00000000000000011001101001010011" ;
			-- 1.843750 => 0.399437
			when "11011000" => x_beta_lut <= "00000000000000011001100100000110" ;
			-- 1.847656 => 0.398170
			when "11011001" => x_beta_lut <= "00000000000000011001011110111010" ;
			-- 1.851563 => 0.396912
			when "11011010" => x_beta_lut <= "00000000000000011001011001110000" ;
			-- 1.855469 => 0.395657
			when "11011011" => x_beta_lut <= "00000000000000011001010100100111" ;
			-- 1.859375 => 0.394413
			when "11011100" => x_beta_lut <= "00000000000000011001001111100001" ;
			-- 1.863281 => 0.393173
			when "11011101" => x_beta_lut <= "00000000000000011001001010011100" ;
			-- 1.867188 => 0.391937
			when "11011110" => x_beta_lut <= "00000000000000011001000101011000" ;
			-- 1.871094 => 0.390713
			when "11011111" => x_beta_lut <= "00000000000000011001000000010111" ;
			-- 1.875000 => 0.389492
			when "11100000" => x_beta_lut <= "00000000000000011000111011010111" ;
			-- 1.878906 => 0.388279
			when "11100001" => x_beta_lut <= "00000000000000011000110110011001" ;
			-- 1.882813 => 0.387070
			when "11100010" => x_beta_lut <= "00000000000000011000110001011100" ;
			-- 1.886719 => 0.385868
			when "11100011" => x_beta_lut <= "00000000000000011000101100100001" ;
			-- 1.890625 => 0.384674
			when "11100100" => x_beta_lut <= "00000000000000011000100111101000" ;
			-- 1.894531 => 0.383484
			when "11100101" => x_beta_lut <= "00000000000000011000100010110000" ;
			-- 1.898438 => 0.382301
			when "11100110" => x_beta_lut <= "00000000000000011000011101111010" ;
			-- 1.902344 => 0.381123
			when "11100111" => x_beta_lut <= "00000000000000011000011001000101" ;
			-- 1.906250 => 0.379951
			when "11101000" => x_beta_lut <= "00000000000000011000010100010010" ;
			-- 1.910156 => 0.378788
			when "11101001" => x_beta_lut <= "00000000000000011000001111100001" ;
			-- 1.914063 => 0.377628
			when "11101010" => x_beta_lut <= "00000000000000011000001010110001" ;
			-- 1.917969 => 0.376476
			when "11101011" => x_beta_lut <= "00000000000000011000000110000011" ;
			-- 1.921875 => 0.375328
			when "11101100" => x_beta_lut <= "00000000000000011000000001010110" ;
			-- 1.925781 => 0.374187
			when "11101101" => x_beta_lut <= "00000000000000010111111100101011" ;
			-- 1.929688 => 0.373051
			when "11101110" => x_beta_lut <= "00000000000000010111111000000001" ;
			-- 1.933594 => 0.371922
			when "11101111" => x_beta_lut <= "00000000000000010111110011011001" ;
			-- 1.937500 => 0.370796
			when "11110000" => x_beta_lut <= "00000000000000010111101110110010" ;
			-- 1.941406 => 0.369678
			when "11110001" => x_beta_lut <= "00000000000000010111101010001101" ;
			-- 1.945313 => 0.368568
			when "11110010" => x_beta_lut <= "00000000000000010111100101101010" ;
			-- 1.949219 => 0.367458
			when "11110011" => x_beta_lut <= "00000000000000010111100001000111" ;
			-- 1.953125 => 0.366356
			when "11110100" => x_beta_lut <= "00000000000000010111011100100110" ;
			-- 1.957031 => 0.365261
			when "11110101" => x_beta_lut <= "00000000000000010111011000000111" ;
			-- 1.960938 => 0.364170
			when "11110110" => x_beta_lut <= "00000000000000010111010011101001" ;
			-- 1.964844 => 0.363083
			when "11110111" => x_beta_lut <= "00000000000000010111001111001100" ;
			-- 1.968750 => 0.362003
			when "11111000" => x_beta_lut <= "00000000000000010111001010110001" ;
			-- 1.972656 => 0.360931
			when "11111001" => x_beta_lut <= "00000000000000010111000110011000" ;
			-- 1.976563 => 0.359859
			when "11111010" => x_beta_lut <= "00000000000000010111000001111111" ;
			-- 1.980469 => 0.358795
			when "11111011" => x_beta_lut <= "00000000000000010110111101101000" ;
			-- 1.984375 => 0.357738
			when "11111100" => x_beta_lut <= "00000000000000010110111001010011" ;
			-- 1.988281 => 0.356682
			when "11111101" => x_beta_lut <= "00000000000000010110110100111110" ;
			-- 1.992188 => 0.355637
			when "11111110" => x_beta_lut <= "00000000000000010110110000101100" ;
			-- 1.996094 => 0.354591
			when "11111111" => x_beta_lut <= "00000000000000010110101100011010" ;
			when others => x_beta_lut <= x"00000000" ;
        end case;
		end if;
    end process;
end architecture; 